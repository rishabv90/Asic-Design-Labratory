// $ID: mg 147$
// File name: flex counter$  
// Author: Rishab Verma     $
// Lab Section: Friday 11 30$
// Description: $




module flex_counter#(
    parameter NUM_CNT_BITS = 4
)
(
    input wire clk,
    input wire n_rst,
    input wire count_enable,
    input wire clear,
    input wire [(NUM_CNT_BITS-1):0] rollover_val,
    output wire rollover_flag,
    output wire [(NUM_CNT_BITS-1):0] count_out
);


reg flagtmp;
reg nextflag;


reg [(NUM_CNT_BITS-1):0] tempnxt;
reg [(NUM_CNT_BITS-1):0] tempcount;


always_ff @ (posedge clk, negedge n_rst)
begin
	if(n_rst == 0)
	begin
	 
		  tempcount <= 0;
	 	  flagtmp <= 1'b0;
	end 
	else 
	begin
	   	tempcount <= tempnxt;
	   	flagtmp <= nextflag;
	end
end
   
always_comb 
begin
      if(clear == 1) 
      begin
	 	tempnxt = 0;
	 	nextflag = 1'b0;
      end 

      else 
      begin
	 if(count_enable == 1) 
	 begin
	 	   tempnxt = tempcount + 1;
	 	   nextflag = 1'b0;

	    if(tempnxt == (rollover_val + 1)) 
	    begin
	 	      tempnxt = 1;
	    end

	    if(tempnxt == rollover_val) 
	    begin
	 	      nextflag = 1'b1;
	    end
	 end 

	else 
	begin
	 	   nextflag = flagtmp;
	 	   tempnxt = tempcount;
	 end 
      end 
   end
   
   assign rollover_flag = flagtmp;
   assign count_out = tempcount;
      

endmodule

/*
`timescale 1ns /100ps

module adder_1bit
(
	input wire a,
	input wire b,
	input wire carry_in,
	
	output reg sum,
	output reg carry_out
);
 
always @ (a,b, carry_in)
   begin
      assert(( a == 1'b1) || (a == 1'b0))
      else $error("Input 'a' of component is not a digital logic value");

      assert((b == 1'b1) || (b == 1'b0))
      else $error("Input 'b' of component is not a digital logic value");

      assert((carry_in == 1'b1) || (carry_in == 1'b0))
      else $error("Input 'carry_in' of component is not a digital logic value");
	
   end



  assign sum = carry_in ^ (a ^ b);
  assign carry_out = ((! carry_in) & b & a) | (carry_in & (b | a));


   
   always @ (a, b, carry_in)
   begin
     #(2) assert (((a+b+carry_in)%2) == sum)
       else $error("Output 's' of first 1 bit adder is not correct");
   end
	

endmodule
`timescale 1ns /100ps

module adder_1bit
(
	input wire a,
	input wire b,
	input wire carry_in,
	
	output reg sum,
	output reg carry_out
);
 
always @ (a,b, carry_in)
   begin
      assert(( a == 1'b1) || (a == 1'b0))
      else $error("Input 'a' of component is not a digital logic value");

      assert((b == 1'b1) || (b == 1'b0))
      else $error("Input 'b' of component is not a digital logic value");

      assert((carry_in == 1'b1) || (carry_in == 1'b0))
      else $error("Input 'carry_in' of component is not a digital logic value");
	
   end



  assign sum = carry_in ^ (a ^ b);
  assign carry_out = ((! carry_in) & b & a) | (carry_in & (b | a));


   
   always @ (a, b, carry_in)
   begin
     #(2) assert (((a+b+carry_in)%2) == sum)
       else $error("Output 's' of first 1 bit adder is not correct");
   end
	

endmodule

*/