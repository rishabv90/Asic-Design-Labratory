
`timescale 1ns / 100ps

module tb_decode
();

	reg tb_clk;
	reg tb_n_rst;
	reg tb_d_plus;
	reg tb_shift_enable;
	reg tb_eop;
	reg tb_d_orig;
	
	localparam CLK_PERIOD = 6;
	localparam CHECK_CLK = 1;
	
	decode DUT (.clk(tb_clk), .n_rst(tb_n_rst), .d_plus(tb_d_plus), .shift_enable(tb_shift_enable), .eop(tb_eop), .d_orig(tb_d_orig) );
	
	
  	always
  	begin : CLK_GEN
   	tb_clk = 1'b0;
    	#(CLK_PERIOD/2);
    	tb_clk = 1'b1;
    	#(CLK_PERIOD/2);
  	end
  	
  initial
  begin
  
	tb_n_rst = 1'b0;
	#(1);
	tb_n_rst = 1'b1;
	
	tb_d_plus = 1'b0; @ (posedge tb_clk);
	tb_shift_enable = 1'b0; @ (posedge tb_clk);
	tb_eop = 1'b0; @ (posedge tb_clk);
	
	#(5);
	tb_d_plus = 1'b1; @ (posedge tb_clk);
	#(5);
	tb_shift_enable = 1'b1; @ (posedge tb_clk); 
	#(1);
	assert(tb_d_orig == 1'b0) 
	begin
		$display("test case 1 passed");
	end 
	else 
	begin
		$error("test case 1 failed");
	end
	#(2);
	tb_shift_enable = 1'b0; @ (posedge tb_clk); 
	
	
	#(5);
	tb_shift_enable = 1'b1; @ (posedge tb_clk); 
	#(1);
	assert(tb_d_orig == 1'b1) 
	begin
		$display("test case 1 passed");
	end 
	else 
	begin
		$error("test case 1 failed");
	end
	#(2);
	tb_shift_enable = 1'b0; @ (posedge tb_clk); 
	
	#(5);
	tb_d_plus = 1'b0; @ (posedge tb_clk);
	#(5);
	tb_shift_enable = 1'b1; @ (posedge tb_clk); 
	#(1);
	assert(tb_d_orig == 1'b0) 
	begin
		$display("test case 1 passed");
	end 
	else 
	begin
		$error("test case 1 failed");
	end
	#(2);
	tb_shift_enable = 1'b0; @ (posedge tb_clk); 
	
  end
  	
endmodule
